magic
tech sky130A
timestamp 1614660232
<< nwell >>
rect -70 100 150 1000
<< nmos >>
rect 0 -130 15 -30
rect 65 -130 80 -30
rect 0 -375 15 -275
<< pmos >>
rect 0 775 15 875
rect 65 775 80 875
rect 0 530 15 630
rect 0 125 15 225
<< ndiff >>
rect -50 -45 0 -30
rect -50 -115 -35 -45
rect -15 -115 0 -45
rect -50 -130 0 -115
rect 15 -45 65 -30
rect 15 -115 30 -45
rect 50 -115 65 -45
rect 15 -130 65 -115
rect 80 -45 130 -30
rect 80 -115 95 -45
rect 115 -115 130 -45
rect 80 -130 130 -115
rect -50 -290 0 -275
rect -50 -360 -35 -290
rect -15 -360 0 -290
rect -50 -375 0 -360
rect 15 -290 60 -275
rect 15 -360 30 -290
rect 50 -360 60 -290
rect 15 -375 60 -360
<< pdiff >>
rect -50 860 0 875
rect -50 790 -35 860
rect -15 790 0 860
rect -50 775 0 790
rect 15 860 65 875
rect 15 790 30 860
rect 50 790 65 860
rect 15 775 65 790
rect 80 860 130 875
rect 80 790 95 860
rect 115 790 130 860
rect 80 775 130 790
rect -50 615 0 630
rect -50 545 -35 615
rect -15 545 0 615
rect -50 530 0 545
rect 15 615 65 630
rect 15 545 30 615
rect 50 545 65 615
rect 15 530 65 545
rect -50 210 0 225
rect -50 140 -35 210
rect -15 140 0 210
rect -50 125 0 140
rect 15 210 65 225
rect 15 140 30 210
rect 50 140 65 210
rect 15 125 65 140
<< ndiffc >>
rect -35 -115 -15 -45
rect 30 -115 50 -45
rect 95 -115 115 -45
rect -35 -360 -15 -290
rect 30 -360 50 -290
<< pdiffc >>
rect -35 790 -15 860
rect 30 790 50 860
rect 95 790 115 860
rect -35 545 -15 615
rect 30 545 50 615
rect -35 140 -15 210
rect 30 140 50 210
<< psubdiff >>
rect 60 -290 110 -275
rect 60 -360 75 -290
rect 95 -360 110 -290
rect 60 -375 110 -360
<< nsubdiff >>
rect -10 955 90 970
rect -10 935 5 955
rect 75 935 90 955
rect -10 920 90 935
<< psubdiffcont >>
rect 75 -360 95 -290
<< nsubdiffcont >>
rect 5 935 75 955
<< poly >>
rect 0 875 15 890
rect 65 875 80 890
rect 0 710 15 775
rect 65 760 80 775
rect 65 745 135 760
rect 0 700 95 710
rect 0 680 10 700
rect 30 695 95 700
rect 30 680 40 695
rect 0 670 40 680
rect 0 630 15 645
rect 0 520 15 530
rect -65 505 15 520
rect -65 320 -50 505
rect 80 480 95 695
rect -25 465 95 480
rect -25 365 -10 465
rect 15 430 55 440
rect 15 410 25 430
rect 45 415 55 430
rect 120 415 135 745
rect 45 410 135 415
rect 15 400 135 410
rect 119 390 160 400
rect 119 369 129 390
rect 148 369 160 390
rect -25 355 95 365
rect 119 360 160 369
rect -25 350 65 355
rect 55 335 65 350
rect 85 335 95 355
rect 55 325 95 335
rect -65 315 15 320
rect -65 305 35 315
rect 0 300 35 305
rect -65 270 -25 280
rect -65 250 -55 270
rect -35 255 -25 270
rect 20 255 35 300
rect -35 250 35 255
rect -65 240 35 250
rect 0 235 35 240
rect 0 225 15 235
rect 0 80 15 125
rect -75 65 15 80
rect -75 -245 -60 65
rect 80 40 95 325
rect 0 25 95 40
rect 0 -30 15 25
rect 120 0 135 360
rect 65 -15 135 0
rect 65 -30 80 -15
rect 0 -145 15 -130
rect 65 -145 80 -130
rect -75 -260 15 -245
rect 0 -275 15 -260
rect 0 -390 15 -375
<< polycont >>
rect 10 680 30 700
rect 25 410 45 430
rect 129 369 148 390
rect 65 335 85 355
rect -55 250 -35 270
<< locali >>
rect -5 955 85 965
rect -5 935 5 955
rect 75 935 85 955
rect -5 925 85 935
rect 30 870 50 925
rect -45 860 -5 870
rect -45 790 -35 860
rect -15 790 -5 860
rect -45 780 -5 790
rect 20 860 60 870
rect 20 790 30 860
rect 50 790 60 860
rect 20 780 60 790
rect 85 860 125 870
rect 85 790 95 860
rect 115 790 125 860
rect 85 780 125 790
rect -25 755 -5 780
rect 105 760 125 780
rect -25 735 80 755
rect 105 740 140 760
rect 0 700 40 710
rect 0 680 10 700
rect 30 680 40 700
rect 0 670 40 680
rect 20 625 40 670
rect 60 670 80 735
rect 60 650 100 670
rect -75 615 -5 625
rect -75 605 -35 615
rect -45 545 -35 605
rect -15 545 -5 615
rect -45 535 -5 545
rect 20 615 60 625
rect 20 545 30 615
rect 50 545 60 615
rect 20 535 60 545
rect 80 510 100 650
rect -25 490 100 510
rect 120 625 140 740
rect 120 605 155 625
rect -25 440 -5 490
rect 120 470 140 605
rect 75 450 140 470
rect -25 430 55 440
rect -25 410 25 430
rect 45 410 55 430
rect -25 400 55 410
rect -25 320 -5 400
rect 75 365 95 450
rect 55 355 95 365
rect 119 390 171 400
rect 119 369 129 390
rect 148 379 171 390
rect 148 369 160 379
rect 119 360 160 369
rect 55 335 65 355
rect 85 335 95 355
rect 55 325 95 335
rect -25 300 35 320
rect 60 305 80 325
rect -65 270 -25 280
rect -65 260 -55 270
rect -75 250 -55 260
rect -35 250 -25 270
rect -75 240 -25 250
rect 17 260 34 300
rect 60 285 140 305
rect 17 240 100 260
rect 80 220 100 240
rect -75 210 -5 220
rect -75 200 -35 210
rect -45 140 -35 200
rect -15 140 -5 210
rect -45 130 -5 140
rect 20 210 100 220
rect 20 140 30 210
rect 50 200 100 210
rect 50 140 60 200
rect 20 130 60 140
rect 80 15 100 200
rect -25 -5 100 15
rect -25 -30 -5 -5
rect -45 -45 -5 -30
rect 120 -35 140 285
rect -45 -115 -35 -45
rect -15 -115 -5 -45
rect -45 -125 -5 -115
rect 20 -45 60 -35
rect 20 -115 30 -45
rect 50 -115 60 -45
rect 20 -125 60 -115
rect 85 -45 140 -35
rect 85 -115 95 -45
rect 115 -65 140 -45
rect 115 -115 125 -65
rect 85 -125 125 -115
rect 20 -200 40 -125
rect -25 -220 40 -200
rect -25 -280 -5 -220
rect -45 -290 -5 -280
rect -45 -360 -35 -290
rect -15 -360 -5 -290
rect -45 -370 -5 -360
rect 20 -290 105 -280
rect 20 -360 30 -290
rect 50 -360 75 -290
rect 95 -360 105 -290
rect 20 -370 105 -360
<< viali >>
rect 5 935 75 955
rect 30 790 50 860
rect 30 -360 50 -290
rect 75 -360 95 -290
<< metal1 >>
rect -75 955 145 1000
rect -75 935 5 955
rect 75 935 145 955
rect -75 875 145 935
rect -76 860 146 875
rect -76 790 30 860
rect 50 790 146 860
rect -76 775 146 790
rect -64 320 146 775
rect -65 300 146 320
rect -64 280 146 300
rect -65 240 146 280
rect -64 123 146 240
rect -68 -290 147 -31
rect -68 -360 30 -290
rect 50 -360 75 -290
rect 95 -360 147 -290
rect -68 -377 147 -360
<< labels >>
rlabel locali -75 615 -75 615 7 D
port 1 w
rlabel locali 155 615 155 615 3 Q
port 3 e
rlabel locali -75 210 -75 210 7 Db
port 2 w
rlabel locali 171 389 171 389 3 Qb
port 4 e
rlabel metal1 -76 825 -76 825 7 VP
port 5 w
rlabel metal1 -68 -326 -68 -326 7 VN
port 6 w
rlabel locali -75 250 -75 250 7 clk
port 7 w
<< end >>
