* SPICE3 file created from CSRL_latch_half_2_top_layout.ext - technology: sky130A

.subckt CSRL_latch_half_2 D Db clk VP VN Q Qb
X0 Q Qb a_1060_880# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X1 Q clk D VN sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X2 VN Q Qb VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X3 Q Qb VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Qb clk Db VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X5 VP clk a_1060_880# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_1060_880# Q Qb VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
.ends


* Top level circuit CSRL_latch_half_2_top_layout

XCSRL_latch_half_2_0 D Db clk VP VN Q Qb CSRL_latch_half_2
.end

