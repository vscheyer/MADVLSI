magic
tech sky130A
timestamp 1614632775
<< locali >>
rect 342 303 372 323
rect -3 263 27 283
rect -3 203 27 223
rect 342 203 372 223
rect -3 18 27 38
<< metal1 >>
rect 7 663 21 763
rect 17 88 31 188
use CSRL_latch_half_2  CSRL_latch_half_2_0 ~/Documents/Mini_Project_2/half_CSRL_2/layout
timestamp 1614632467
transform 1 0 -413 0 1 478
box 410 -480 785 560
<< labels >>
rlabel metal1 7 733 7 733 7 VP
rlabel locali -3 273 -3 273 7 Db
rlabel locali -3 213 -3 213 7 D
rlabel metal1 17 138 17 138 7 VN
rlabel locali -3 28 -3 28 7 clk
rlabel locali 372 313 372 313 3 Q
rlabel locali 372 213 372 213 3 Qb
<< end >>
