magic
tech sky130A
timestamp 1613685484
<< nwell >>
rect -120 135 290 275
<< nmos >>
rect 0 0 15 100
rect 205 0 220 100
<< pmos >>
rect 0 155 15 255
rect 205 155 220 255
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 155 85 205 100
rect 155 15 170 85
rect 190 15 205 85
rect 155 0 205 15
rect 220 85 270 100
rect 220 15 235 85
rect 255 15 270 85
rect 220 0 270 15
<< pdiff >>
rect -50 240 0 255
rect -50 170 -35 240
rect -15 170 0 240
rect -50 155 0 170
rect 15 240 65 255
rect 15 170 30 240
rect 50 170 65 240
rect 15 155 65 170
rect 155 240 205 255
rect 155 170 170 240
rect 190 170 205 240
rect 155 155 205 170
rect 220 240 270 255
rect 220 170 235 240
rect 255 170 270 240
rect 220 155 270 170
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
rect 170 15 190 85
rect 235 15 255 85
<< pdiffc >>
rect -35 170 -15 240
rect 30 170 50 240
rect 170 170 190 240
rect 235 170 255 240
<< psubdiff >>
rect -100 85 -50 100
rect -100 15 -85 85
rect -65 15 -50 85
rect -100 0 -50 15
<< nsubdiff >>
rect -100 240 -50 255
rect -100 170 -85 240
rect -65 170 -50 240
rect -100 155 -50 170
rect 105 240 155 255
rect 105 170 120 240
rect 140 170 155 240
rect 105 155 155 170
<< psubdiffcont >>
rect -85 15 -65 85
<< nsubdiffcont >>
rect -85 170 -65 240
rect 120 170 140 240
<< poly >>
rect 0 255 15 270
rect 205 255 220 270
rect 0 100 15 155
rect 205 100 220 155
rect 0 -15 15 0
rect 205 -15 220 0
rect -25 -25 15 -15
rect -25 -45 -15 -25
rect 5 -45 15 -25
rect -25 -55 15 -45
rect 180 -25 220 -15
rect 180 -45 190 -25
rect 210 -45 220 -25
rect 180 -55 220 -45
<< polycont >>
rect -15 -45 5 -25
rect 190 -45 210 -25
<< locali >>
rect -95 240 -5 250
rect -95 170 -85 240
rect -65 170 -35 240
rect -15 170 -5 240
rect -95 160 -5 170
rect 20 240 60 250
rect 20 170 30 240
rect 50 170 60 240
rect 20 160 60 170
rect 110 240 200 250
rect 110 170 120 240
rect 140 170 170 240
rect 190 170 200 240
rect 110 160 200 170
rect 225 240 265 250
rect 225 170 235 240
rect 255 170 265 240
rect 225 160 265 170
rect 40 134 60 160
rect 245 134 265 160
rect 40 114 292 134
rect 245 95 265 114
rect -95 85 -5 95
rect -95 15 -85 85
rect -65 15 -35 85
rect -15 15 -5 85
rect -95 5 -5 15
rect 20 85 60 95
rect 20 15 30 85
rect 50 25 60 85
rect 110 85 200 95
rect 110 25 170 85
rect 50 15 170 25
rect 190 15 200 85
rect 20 5 200 15
rect 225 85 265 95
rect 225 15 235 85
rect 255 15 265 85
rect 225 5 265 15
rect -120 -25 15 -15
rect -120 -35 -15 -25
rect -25 -45 -15 -35
rect 5 -45 15 -25
rect 85 -25 220 -15
rect 85 -35 190 -25
rect -25 -55 15 -45
rect 180 -45 190 -35
rect 210 -45 220 -25
rect 180 -55 220 -45
<< viali >>
rect -85 170 -65 240
rect -35 170 -15 240
rect 120 170 140 240
rect 170 170 190 240
rect -85 15 -65 85
rect -35 15 -15 85
<< metal1 >>
rect -120 240 290 250
rect -120 170 -85 240
rect -65 170 -35 240
rect -15 170 120 240
rect 140 170 170 240
rect 190 170 290 240
rect -120 160 290 170
rect -120 85 290 95
rect -120 15 -85 85
rect -65 15 -35 85
rect -15 15 290 85
rect -120 5 290 15
<< labels >>
rlabel locali -120 -25 -120 -25 7 A
port 1 w
rlabel metal1 -120 205 -120 205 7 VP
port 3 w
rlabel metal1 -120 50 -120 50 7 VN
port 4 w
rlabel locali 85 -25 85 -25 7 B
port 2 w
rlabel locali 292 124 292 124 3 Y
port 5 e
<< end >>
