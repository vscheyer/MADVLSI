magic
tech sky130A
timestamp 1614710634
<< nwell >>
rect -75 986 400 1000
rect -75 765 401 986
rect -75 510 400 765
rect -75 100 150 510
<< nmos >>
rect 240 125 255 225
rect 0 -230 15 -130
rect 65 -230 80 -130
rect 240 -230 255 -130
rect 0 -475 15 -375
rect 240 -475 255 -375
rect 305 -475 320 -375
<< pmos >>
rect 0 775 15 875
rect 65 775 80 875
rect 305 775 320 875
rect 0 530 15 630
rect 0 125 15 225
rect 240 530 255 630
rect 305 530 320 630
<< ndiff >>
rect 190 210 240 225
rect 190 140 205 210
rect 225 140 240 210
rect 190 125 240 140
rect 255 210 305 225
rect 255 140 270 210
rect 290 140 305 210
rect 255 125 305 140
rect -50 -145 0 -130
rect -50 -215 -35 -145
rect -15 -215 0 -145
rect -50 -230 0 -215
rect 15 -145 65 -130
rect 15 -215 30 -145
rect 50 -215 65 -145
rect 15 -230 65 -215
rect 80 -145 130 -130
rect 80 -215 95 -145
rect 115 -215 130 -145
rect 80 -230 130 -215
rect 190 -145 240 -130
rect 190 -215 205 -145
rect 225 -215 240 -145
rect 190 -230 240 -215
rect 255 -145 305 -130
rect 255 -215 270 -145
rect 290 -215 305 -145
rect 255 -230 305 -215
rect -50 -390 0 -375
rect -50 -460 -35 -390
rect -15 -460 0 -390
rect -50 -475 0 -460
rect 15 -390 60 -375
rect 15 -460 30 -390
rect 50 -460 60 -390
rect 15 -475 60 -460
rect 190 -390 240 -375
rect 190 -460 205 -390
rect 225 -460 240 -390
rect 190 -475 240 -460
rect 255 -390 305 -375
rect 255 -460 270 -390
rect 290 -460 305 -390
rect 255 -475 305 -460
rect 320 -390 370 -375
rect 320 -460 335 -390
rect 355 -460 370 -390
rect 320 -475 370 -460
<< pdiff >>
rect -50 860 0 875
rect -50 790 -35 860
rect -15 790 0 860
rect -50 775 0 790
rect 15 860 65 875
rect 15 790 30 860
rect 50 790 65 860
rect 15 775 65 790
rect 80 860 130 875
rect 80 790 95 860
rect 115 790 130 860
rect 80 775 130 790
rect 255 860 305 875
rect 255 790 270 860
rect 290 790 305 860
rect 255 775 305 790
rect 320 860 370 875
rect 320 790 335 860
rect 355 790 370 860
rect 320 775 370 790
rect -50 615 0 630
rect -50 545 -35 615
rect -15 545 0 615
rect -50 530 0 545
rect 15 615 65 630
rect 15 545 30 615
rect 50 545 65 615
rect 15 530 65 545
rect -50 210 0 225
rect -50 140 -35 210
rect -15 140 0 210
rect -50 125 0 140
rect 15 210 65 225
rect 15 140 30 210
rect 50 140 65 210
rect 15 125 65 140
rect 190 615 240 630
rect 190 545 205 615
rect 225 545 240 615
rect 190 530 240 545
rect 255 615 305 630
rect 255 545 270 615
rect 290 545 305 615
rect 255 530 305 545
rect 320 615 370 630
rect 320 545 335 615
rect 355 545 370 615
rect 320 530 370 545
<< ndiffc >>
rect 205 140 225 210
rect 270 140 290 210
rect -35 -215 -15 -145
rect 30 -215 50 -145
rect 95 -215 115 -145
rect 205 -215 225 -145
rect 270 -215 290 -145
rect -35 -460 -15 -390
rect 30 -460 50 -390
rect 205 -460 225 -390
rect 270 -460 290 -390
rect 335 -460 355 -390
<< pdiffc >>
rect -35 790 -15 860
rect 30 790 50 860
rect 95 790 115 860
rect 270 790 290 860
rect 335 790 355 860
rect -35 545 -15 615
rect 30 545 50 615
rect -35 140 -15 210
rect 30 140 50 210
rect 205 545 225 615
rect 270 545 290 615
rect 335 545 355 615
<< psubdiff >>
rect 60 -390 110 -375
rect 60 -460 75 -390
rect 95 -460 110 -390
rect 60 -475 110 -460
rect 230 -520 330 -505
rect 230 -540 245 -520
rect 315 -540 330 -520
rect 230 -555 330 -540
<< nsubdiff >>
rect -10 955 90 970
rect -10 935 5 955
rect 75 935 90 955
rect -10 920 90 935
rect 205 860 255 875
rect 205 790 220 860
rect 240 790 255 860
rect 205 775 255 790
<< psubdiffcont >>
rect 75 -460 95 -390
rect 245 -540 315 -520
<< nsubdiffcont >>
rect 5 935 75 955
rect 220 790 240 860
<< poly >>
rect 0 875 15 890
rect 65 875 80 890
rect 305 875 320 890
rect 0 720 15 775
rect 65 760 80 775
rect 65 745 140 760
rect 0 710 40 720
rect -65 685 -25 695
rect -65 665 -55 685
rect -35 665 -25 685
rect 0 690 10 710
rect 30 695 95 710
rect 30 690 40 695
rect 0 680 40 690
rect -65 655 -25 665
rect -40 640 15 655
rect 0 630 15 640
rect 0 520 15 530
rect -65 505 15 520
rect -65 320 -50 505
rect 80 480 95 695
rect -25 465 95 480
rect -25 365 -10 465
rect 15 430 55 440
rect 15 410 25 430
rect 45 415 55 430
rect 125 415 140 745
rect 305 740 320 775
rect 45 410 140 415
rect 15 400 140 410
rect -25 355 95 365
rect -25 350 65 355
rect 55 335 65 350
rect 85 335 95 355
rect 55 325 95 335
rect -65 315 15 320
rect -65 305 35 315
rect 0 300 35 305
rect 20 255 35 300
rect 0 235 35 255
rect 0 225 15 235
rect 0 80 15 125
rect -75 65 15 80
rect -75 -345 -60 65
rect 80 -55 95 325
rect 0 -70 95 -55
rect 0 -130 15 -70
rect 125 -75 140 400
rect 165 725 320 740
rect 165 250 180 725
rect 305 695 320 725
rect 305 685 380 695
rect 305 680 350 685
rect 340 665 350 680
rect 370 665 380 685
rect 340 655 380 665
rect 240 630 255 645
rect 305 630 320 645
rect 240 520 255 530
rect 205 505 255 520
rect 305 520 320 530
rect 305 505 375 520
rect 205 415 220 505
rect 245 470 285 480
rect 245 450 255 470
rect 275 455 285 470
rect 360 455 375 505
rect 275 450 375 455
rect 245 440 375 450
rect 205 405 280 415
rect 205 400 250 405
rect 240 385 250 400
rect 270 385 280 405
rect 240 375 280 385
rect 240 315 255 375
rect 240 305 335 315
rect 240 300 265 305
rect 255 285 265 300
rect 285 300 335 305
rect 285 285 295 300
rect 255 275 295 285
rect 165 235 255 250
rect 240 225 255 235
rect 240 115 255 125
rect 320 115 335 300
rect 195 100 255 115
rect 280 100 335 115
rect 125 -85 165 -75
rect 125 -100 135 -85
rect 65 -105 135 -100
rect 155 -105 165 -85
rect 65 -115 165 -105
rect 195 -105 210 100
rect 280 -105 295 100
rect 360 20 375 440
rect 335 10 375 20
rect 335 -10 345 10
rect 365 -10 375 10
rect 335 -20 375 -10
rect 65 -130 80 -115
rect 195 -120 255 -105
rect 280 -120 335 -105
rect 240 -130 255 -120
rect 0 -245 15 -230
rect 65 -245 80 -230
rect 240 -270 255 -230
rect 145 -285 255 -270
rect 145 -345 160 -285
rect 320 -310 335 -120
rect -75 -360 160 -345
rect 240 -325 335 -310
rect 0 -375 15 -360
rect 240 -375 255 -325
rect 360 -350 375 -20
rect 305 -365 375 -350
rect 305 -375 320 -365
rect 0 -490 15 -475
rect 240 -490 255 -475
rect 305 -490 320 -475
<< polycont >>
rect -55 665 -35 685
rect 10 690 30 710
rect 25 410 45 430
rect 65 335 85 355
rect 350 665 370 685
rect 255 450 275 470
rect 250 385 270 405
rect 265 285 285 305
rect 135 -105 155 -85
rect 345 -10 365 10
<< locali >>
rect -5 955 85 965
rect -5 935 5 955
rect 75 935 85 955
rect -5 925 85 935
rect 30 870 50 925
rect -45 860 -5 870
rect -45 790 -35 860
rect -15 790 -5 860
rect -45 780 -5 790
rect 20 860 60 870
rect 20 790 30 860
rect 50 790 60 860
rect 20 780 60 790
rect 85 860 125 870
rect 85 790 95 860
rect 115 790 125 860
rect 85 780 125 790
rect 210 860 300 870
rect 210 790 220 860
rect 240 790 270 860
rect 290 790 300 860
rect 210 780 300 790
rect 325 860 365 870
rect 325 790 335 860
rect 355 790 365 860
rect 325 780 365 790
rect -25 760 -5 780
rect 105 760 125 780
rect -25 740 80 760
rect 105 740 140 760
rect 325 745 345 780
rect 0 710 40 720
rect -65 685 -25 695
rect -65 675 -55 685
rect -75 665 -55 675
rect -35 665 -25 685
rect 0 690 10 710
rect 30 690 40 710
rect 0 680 40 690
rect -75 655 -25 665
rect 20 625 40 680
rect 60 670 80 740
rect 60 650 100 670
rect -75 615 -5 625
rect -75 605 -35 615
rect -45 545 -35 605
rect -15 545 -5 615
rect -45 535 -5 545
rect 20 615 60 625
rect 20 545 30 615
rect 50 545 60 615
rect 20 535 60 545
rect 80 510 100 650
rect -25 490 100 510
rect -25 440 -5 490
rect 120 470 140 740
rect 280 725 345 745
rect 280 625 300 725
rect 340 685 380 695
rect 340 665 350 685
rect 370 675 380 685
rect 370 665 400 675
rect 340 655 400 665
rect 195 615 235 625
rect 195 545 205 615
rect 225 545 235 615
rect 195 535 235 545
rect 260 615 300 625
rect 260 545 270 615
rect 290 545 300 615
rect 260 535 300 545
rect 325 615 400 625
rect 325 545 335 615
rect 355 605 400 615
rect 355 545 365 605
rect 325 535 365 545
rect 75 450 140 470
rect 215 480 235 535
rect 325 510 345 535
rect 315 495 345 510
rect 215 470 285 480
rect 215 460 255 470
rect 195 450 255 460
rect 275 450 285 470
rect -25 430 55 440
rect -25 410 25 430
rect 45 410 55 430
rect -25 400 55 410
rect -25 320 -5 400
rect 75 365 95 450
rect 55 355 95 365
rect 55 335 65 355
rect 85 335 95 355
rect 195 440 285 450
rect 195 355 215 440
rect 240 405 280 415
rect 240 385 250 405
rect 270 395 280 405
rect 315 395 335 495
rect 270 385 380 395
rect 240 375 380 385
rect 195 335 340 355
rect 55 325 95 335
rect -25 300 35 320
rect 60 305 80 325
rect 255 305 295 315
rect 17 260 34 300
rect 60 285 140 305
rect 17 240 100 260
rect 80 220 100 240
rect -45 210 -5 220
rect -45 140 -35 210
rect -15 140 -5 210
rect -45 130 -5 140
rect 20 210 100 220
rect 20 140 30 210
rect 50 200 100 210
rect 50 140 60 200
rect 20 130 60 140
rect -45 10 -25 130
rect -85 -10 -25 10
rect 80 5 100 200
rect 45 -15 100 5
rect 120 185 140 285
rect 255 285 265 305
rect 285 285 295 305
rect 255 275 295 285
rect 275 220 295 275
rect 195 210 235 220
rect 195 185 205 210
rect 120 160 205 185
rect 45 -95 65 -15
rect 120 -35 140 160
rect 195 140 205 160
rect 225 140 235 210
rect 195 130 235 140
rect 260 210 300 220
rect 260 140 270 210
rect 290 140 300 210
rect 260 130 300 140
rect 320 110 340 335
rect -25 -115 65 -95
rect 85 -55 140 -35
rect 245 90 340 110
rect -25 -130 -5 -115
rect -45 -145 -5 -130
rect 85 -135 105 -55
rect 125 -85 165 -75
rect 125 -105 135 -85
rect 155 -95 165 -85
rect 245 -95 265 90
rect 360 70 380 375
rect 285 50 380 70
rect 285 -55 305 50
rect 335 10 375 20
rect 335 -10 345 10
rect 365 -10 390 10
rect 335 -20 375 -10
rect 360 -55 380 -50
rect 285 -75 380 -55
rect 155 -105 215 -95
rect 125 -115 215 -105
rect 245 -115 340 -95
rect 195 -135 215 -115
rect 320 -135 340 -115
rect -45 -215 -35 -145
rect -15 -215 -5 -145
rect -45 -225 -5 -215
rect 20 -145 60 -135
rect 20 -215 30 -145
rect 50 -215 60 -145
rect 20 -225 60 -215
rect 85 -145 125 -135
rect 85 -215 95 -145
rect 115 -215 125 -145
rect 85 -225 125 -215
rect 195 -145 235 -135
rect 195 -215 205 -145
rect 225 -215 235 -145
rect 195 -225 235 -215
rect 260 -145 340 -135
rect 260 -215 270 -145
rect 290 -155 340 -145
rect 290 -215 300 -155
rect 260 -225 300 -215
rect 20 -300 40 -225
rect -25 -320 40 -300
rect -25 -380 -5 -320
rect 320 -340 340 -155
rect 215 -360 340 -340
rect 215 -380 235 -360
rect 360 -380 380 -75
rect -45 -390 -5 -380
rect -45 -460 -35 -390
rect -15 -460 -5 -390
rect -45 -470 -5 -460
rect 20 -390 105 -380
rect 20 -460 30 -390
rect 50 -460 75 -390
rect 95 -460 105 -390
rect 20 -470 105 -460
rect 195 -390 235 -380
rect 195 -460 205 -390
rect 225 -460 235 -390
rect 195 -470 235 -460
rect 260 -390 300 -380
rect 260 -460 270 -390
rect 290 -460 300 -390
rect 260 -470 300 -460
rect 325 -390 380 -380
rect 325 -460 335 -390
rect 355 -410 380 -390
rect 355 -460 365 -410
rect 325 -470 365 -460
rect 270 -510 290 -470
rect 235 -520 325 -510
rect 235 -540 245 -520
rect 315 -540 325 -520
rect 235 -550 325 -540
<< viali >>
rect 5 935 75 955
rect 30 790 50 860
rect 220 790 240 860
rect 270 790 290 860
rect 30 -460 50 -390
rect 75 -460 95 -390
rect 270 -460 290 -390
rect 245 -540 315 -520
<< metal1 >>
rect -75 985 -59 986
rect 385 985 401 986
rect -75 955 401 985
rect -75 935 5 955
rect 75 935 401 955
rect -75 860 401 935
rect -75 790 30 860
rect 50 790 220 860
rect 240 790 270 860
rect 290 790 401 860
rect -75 765 401 790
rect -85 -390 390 -360
rect -85 -460 30 -390
rect 50 -460 75 -390
rect 95 -460 270 -390
rect 290 -460 390 -390
rect -85 -520 390 -460
rect -85 -540 245 -520
rect 315 -540 390 -520
rect -85 -570 390 -540
<< labels >>
rlabel locali -75 615 -75 615 7 D
port 1 w
rlabel locali -85 0 -85 0 7 Db
port 3 w
rlabel locali 390 0 390 0 3 Qb
port 9 e
rlabel locali -75 665 -75 665 7 clk
port 4 w
rlabel locali 400 615 400 615 3 Q
port 10 e
rlabel metal1 -75 825 -75 825 7 VP
port 11 w
rlabel metal1 -85 -425 -85 -425 7 VN
port 12 w
<< end >>
