magic
tech sky130A
timestamp 1614575639
<< nwell >>
rect -90 185 230 540
<< nmos >>
rect 0 -25 15 75
rect 65 -25 80 75
rect 0 -220 15 -120
<< pmos >>
rect 0 415 15 515
rect 145 415 160 515
rect 0 205 15 305
rect 65 205 80 305
<< ndiff >>
rect -50 60 0 75
rect -50 -10 -35 60
rect -15 -10 0 60
rect -50 -25 0 -10
rect 15 60 65 75
rect 15 -10 30 60
rect 50 -10 65 60
rect 15 -25 65 -10
rect 80 60 130 75
rect 80 -10 95 60
rect 115 -10 130 60
rect 80 -25 130 -10
rect -50 -135 0 -120
rect -50 -205 -35 -135
rect -15 -205 0 -135
rect -50 -220 0 -205
rect 15 -135 65 -120
rect 15 -205 30 -135
rect 50 -205 65 -135
rect 15 -220 65 -205
<< pdiff >>
rect -50 500 0 515
rect -50 430 -35 500
rect -15 430 0 500
rect -50 415 0 430
rect 15 500 65 515
rect 15 430 30 500
rect 50 430 65 500
rect 15 415 65 430
rect 95 500 145 515
rect 95 430 110 500
rect 130 430 145 500
rect 95 415 145 430
rect 160 500 210 515
rect 160 430 175 500
rect 195 430 210 500
rect 160 415 210 430
rect -50 290 0 305
rect -50 220 -35 290
rect -15 220 0 290
rect -50 205 0 220
rect 15 290 65 305
rect 15 220 30 290
rect 50 220 65 290
rect 15 205 65 220
rect 80 290 130 305
rect 80 220 95 290
rect 115 220 130 290
rect 80 205 130 220
<< ndiffc >>
rect -35 -10 -15 60
rect 30 -10 50 60
rect 95 -10 115 60
rect -35 -205 -15 -135
rect 30 -205 50 -135
<< pdiffc >>
rect -35 430 -15 500
rect 30 430 50 500
rect 110 430 130 500
rect 175 430 195 500
rect -35 220 -15 290
rect 30 220 50 290
rect 95 220 115 290
<< psubdiff >>
rect 140 -70 190 -55
rect 140 -140 155 -70
rect 175 -140 190 -70
rect 140 -155 190 -140
<< nsubdiff >>
rect 157 290 207 305
rect 157 220 172 290
rect 192 220 207 290
rect 157 205 207 220
<< psubdiffcont >>
rect 155 -140 175 -70
<< nsubdiffcont >>
rect 172 220 192 290
<< poly >>
rect 0 515 15 530
rect 145 515 160 530
rect 0 400 15 415
rect 145 400 160 415
rect -65 390 160 400
rect -65 370 -55 390
rect -35 385 160 390
rect -35 370 -25 385
rect -65 360 -25 370
rect 0 350 145 360
rect 0 345 115 350
rect 0 305 15 345
rect 105 330 115 345
rect 135 330 145 350
rect 105 320 145 330
rect 65 305 80 320
rect 0 130 15 205
rect 65 190 80 205
rect 45 180 85 190
rect 45 160 55 180
rect 75 160 85 180
rect 45 150 85 160
rect 155 165 195 175
rect 155 150 165 165
rect 65 145 165 150
rect 185 145 195 165
rect 65 135 195 145
rect -5 120 35 130
rect -5 100 5 120
rect 25 100 35 120
rect -5 90 35 100
rect 0 75 15 90
rect 65 75 80 135
rect 0 -40 15 -25
rect 65 -40 80 -25
rect -25 -75 15 -65
rect -25 -95 -15 -75
rect 5 -95 15 -75
rect -25 -105 15 -95
rect 0 -120 15 -105
rect 0 -235 15 -220
<< polycont >>
rect -55 370 -35 390
rect 115 330 135 350
rect 55 160 75 180
rect 165 145 185 165
rect 5 100 25 120
rect -15 -95 5 -75
<< locali >>
rect -45 510 -25 555
rect 100 510 120 555
rect -45 500 -5 510
rect -45 430 -35 500
rect -15 430 -5 500
rect -45 420 -5 430
rect 20 500 60 510
rect 20 430 30 500
rect 50 430 60 500
rect 20 420 60 430
rect 100 500 140 510
rect 100 430 110 500
rect 130 430 140 500
rect 100 420 140 430
rect 165 500 205 510
rect 165 430 175 500
rect 195 430 205 500
rect 165 420 205 430
rect -65 390 -25 400
rect -65 380 -55 390
rect -85 370 -55 380
rect -35 370 -25 390
rect -85 360 -25 370
rect -85 -65 -65 360
rect 40 340 60 420
rect 185 360 205 420
rect -45 320 60 340
rect 105 350 205 360
rect 105 330 115 350
rect 135 340 205 350
rect 135 330 145 340
rect 105 320 145 330
rect -45 300 -25 320
rect -45 290 -5 300
rect -45 220 -35 290
rect -15 220 -5 290
rect -45 210 -5 220
rect 20 290 60 300
rect 20 220 30 290
rect 50 220 60 290
rect 20 210 60 220
rect 85 290 130 300
rect 85 220 95 290
rect 115 220 130 290
rect 85 210 130 220
rect 157 290 202 300
rect 157 220 172 290
rect 192 220 202 290
rect 157 210 202 220
rect -45 190 -25 210
rect -45 180 85 190
rect -45 170 55 180
rect -45 70 -25 170
rect 45 160 55 170
rect 75 160 85 180
rect 45 150 85 160
rect -5 120 35 130
rect -5 100 5 120
rect 25 110 35 120
rect 105 110 125 210
rect 155 165 195 175
rect 155 145 165 165
rect 185 155 195 165
rect 185 145 230 155
rect 155 135 230 145
rect 25 100 230 110
rect -5 90 230 100
rect 105 70 125 90
rect -45 60 -5 70
rect -45 -10 -35 60
rect -15 -10 -5 60
rect -45 -20 -5 -10
rect 20 60 60 70
rect 20 -10 30 60
rect 50 -10 60 60
rect 20 -20 60 -10
rect 85 60 130 70
rect 85 -10 95 60
rect 115 -10 130 60
rect 85 -20 130 -10
rect -85 -75 15 -65
rect -85 -85 -15 -75
rect -25 -95 -15 -85
rect 5 -95 15 -75
rect -25 -105 15 -95
rect 40 -125 60 -20
rect -45 -135 -5 -125
rect -45 -205 -35 -135
rect -15 -205 -5 -135
rect -45 -215 -5 -205
rect 20 -135 60 -125
rect 20 -205 30 -135
rect 50 -205 60 -135
rect 140 -70 185 -60
rect 140 -140 155 -70
rect 175 -140 185 -70
rect 140 -150 185 -140
rect 20 -215 60 -205
<< viali >>
rect 30 220 50 290
rect 172 220 192 290
rect -35 -205 -15 -135
rect 155 -140 175 -70
<< metal1 >>
rect -65 290 225 515
rect -65 220 30 290
rect 50 220 172 290
rect 192 220 225 290
rect -65 205 225 220
rect -65 -70 195 75
rect -65 -135 155 -70
rect -65 -205 -35 -135
rect -15 -140 155 -135
rect 175 -140 195 -70
rect -15 -205 195 -140
rect -65 -220 195 -205
<< labels >>
rlabel locali -35 555 -35 555 1 Db
port 2 n
rlabel locali 110 555 110 555 1 D
port 1 n
rlabel locali -85 -75 -85 -75 7 clk
port 5 w
rlabel locali 230 100 230 100 3 Q
port 3 e
rlabel locali 230 145 230 145 3 Qb
port 4 e
rlabel metal1 -65 465 -65 465 7 VP
port 6 w
rlabel metal1 -65 -170 -65 -170 7 VN
port 7 w
<< end >>
