magic
tech sky130A
timestamp 1614632467
<< nwell >>
rect 430 185 730 560
<< nmos >>
rect 580 -130 595 -30
rect 645 -130 660 -30
rect 500 -390 515 -290
rect 645 -390 660 -290
<< pmos >>
rect 580 440 595 540
rect 580 205 595 305
rect 645 205 660 305
<< ndiff >>
rect 530 -45 580 -30
rect 530 -115 545 -45
rect 565 -115 580 -45
rect 530 -130 580 -115
rect 595 -45 645 -30
rect 595 -115 610 -45
rect 630 -115 645 -45
rect 595 -130 645 -115
rect 660 -45 710 -30
rect 660 -115 675 -45
rect 695 -115 710 -45
rect 660 -130 710 -115
rect 450 -305 500 -290
rect 450 -375 465 -305
rect 485 -375 500 -305
rect 450 -390 500 -375
rect 515 -305 565 -290
rect 515 -375 530 -305
rect 550 -375 565 -305
rect 515 -390 565 -375
rect 595 -305 645 -290
rect 595 -375 610 -305
rect 630 -375 645 -305
rect 595 -390 645 -375
rect 660 -305 710 -290
rect 660 -375 675 -305
rect 695 -375 710 -305
rect 660 -390 710 -375
<< pdiff >>
rect 530 525 580 540
rect 530 455 545 525
rect 565 455 580 525
rect 530 440 580 455
rect 595 525 645 540
rect 595 455 610 525
rect 630 455 645 525
rect 595 440 645 455
rect 530 290 580 305
rect 530 220 545 290
rect 565 220 580 290
rect 530 205 580 220
rect 595 290 645 305
rect 595 220 610 290
rect 630 220 645 290
rect 595 205 645 220
rect 660 290 710 305
rect 660 220 675 290
rect 695 220 710 290
rect 660 205 710 220
<< ndiffc >>
rect 545 -115 565 -45
rect 610 -115 630 -45
rect 675 -115 695 -45
rect 465 -375 485 -305
rect 530 -375 550 -305
rect 610 -375 630 -305
rect 675 -375 695 -305
<< pdiffc >>
rect 545 455 565 525
rect 610 455 630 525
rect 545 220 565 290
rect 610 220 630 290
rect 675 220 695 290
<< psubdiff >>
rect 570 35 670 50
rect 570 15 585 35
rect 655 15 670 35
rect 570 0 670 15
<< nsubdiff >>
rect 645 525 694 540
rect 645 455 660 525
rect 680 455 694 525
rect 645 440 694 455
<< psubdiffcont >>
rect 585 15 655 35
<< nsubdiffcont >>
rect 660 455 680 525
<< poly >>
rect 580 540 595 555
rect 580 415 595 440
rect 500 400 595 415
rect 500 -290 515 400
rect 580 305 595 320
rect 645 305 660 320
rect 580 125 595 205
rect 645 190 660 205
rect 620 180 660 190
rect 620 160 630 180
rect 650 160 660 180
rect 620 150 660 160
rect 580 115 620 125
rect 580 100 590 115
rect 540 95 590 100
rect 610 95 620 115
rect 540 85 620 95
rect 645 100 660 150
rect 645 85 700 100
rect 540 -5 555 85
rect 685 -5 700 85
rect 540 -20 595 -5
rect 580 -30 595 -20
rect 645 -20 700 -5
rect 645 -30 660 -20
rect 580 -140 595 -130
rect 540 -155 595 -140
rect 540 -235 555 -155
rect 645 -195 660 -130
rect 645 -205 725 -195
rect 645 -210 695 -205
rect 685 -225 695 -210
rect 715 -225 725 -205
rect 685 -235 725 -225
rect 540 -245 580 -235
rect 540 -265 550 -245
rect 570 -265 580 -245
rect 540 -275 580 -265
rect 645 -290 660 -275
rect 500 -400 515 -390
rect 645 -400 660 -390
rect 500 -415 660 -400
rect 645 -440 660 -415
rect 620 -450 660 -440
rect 620 -470 630 -450
rect 650 -470 660 -450
rect 620 -480 660 -470
<< polycont >>
rect 630 160 650 180
rect 590 95 610 115
rect 695 -225 715 -205
rect 550 -265 570 -245
rect 630 -470 650 -450
<< locali >>
rect 535 525 575 535
rect 535 455 545 525
rect 565 455 575 525
rect 535 445 575 455
rect 600 525 690 535
rect 600 455 610 525
rect 630 455 660 525
rect 680 455 690 525
rect 600 445 690 455
rect 555 340 575 445
rect 555 320 620 340
rect 600 300 620 320
rect 535 290 575 300
rect 535 220 545 290
rect 565 220 575 290
rect 535 210 575 220
rect 600 290 640 300
rect 600 220 610 290
rect 630 220 640 290
rect 600 210 640 220
rect 665 290 705 300
rect 665 220 675 290
rect 695 220 705 290
rect 665 210 705 220
rect 535 190 555 210
rect 535 180 660 190
rect 535 170 630 180
rect 535 145 555 170
rect 620 160 630 170
rect 650 160 660 180
rect 620 150 660 160
rect 500 125 555 145
rect 500 5 520 125
rect 580 115 620 125
rect 580 95 590 115
rect 610 105 620 115
rect 685 105 705 210
rect 610 95 705 105
rect 580 85 705 95
rect 575 35 665 45
rect 575 15 585 35
rect 655 15 665 35
rect 575 5 665 15
rect 500 -15 555 5
rect 535 -35 555 -15
rect 609 -35 630 5
rect 685 -35 705 85
rect 530 -45 575 -35
rect 530 -115 545 -45
rect 565 -115 575 -45
rect 530 -125 575 -115
rect 600 -45 640 -35
rect 600 -115 610 -45
rect 630 -115 640 -45
rect 600 -125 640 -115
rect 665 -45 705 -35
rect 665 -115 675 -45
rect 695 -115 705 -45
rect 665 -125 705 -115
rect 555 -155 575 -125
rect 685 -155 705 -125
rect 555 -175 660 -155
rect 685 -175 785 -155
rect 410 -215 620 -195
rect 540 -245 580 -235
rect 410 -275 475 -255
rect 455 -295 475 -275
rect 540 -265 550 -245
rect 570 -265 580 -245
rect 540 -275 580 -265
rect 540 -295 560 -275
rect 455 -305 495 -295
rect 455 -375 465 -305
rect 485 -375 495 -305
rect 455 -385 495 -375
rect 520 -305 560 -295
rect 520 -375 530 -305
rect 550 -375 560 -305
rect 520 -385 560 -375
rect 600 -295 620 -215
rect 640 -255 660 -175
rect 685 -205 725 -195
rect 685 -225 695 -205
rect 715 -225 725 -205
rect 685 -235 725 -225
rect 705 -255 725 -235
rect 640 -275 685 -255
rect 705 -275 785 -255
rect 665 -295 685 -275
rect 600 -305 640 -295
rect 600 -375 610 -305
rect 630 -375 640 -305
rect 600 -385 640 -375
rect 665 -305 705 -295
rect 665 -375 675 -305
rect 695 -375 705 -305
rect 665 -385 705 -375
rect 410 -450 660 -440
rect 410 -460 630 -450
rect 620 -470 630 -460
rect 650 -470 660 -450
rect 620 -480 660 -470
<< viali >>
rect 610 455 630 525
rect 660 455 680 525
rect 585 15 655 35
rect 610 -115 630 -45
<< metal1 >>
rect 420 525 730 550
rect 420 455 610 525
rect 630 455 660 525
rect 680 455 730 525
rect 420 185 730 455
rect 430 35 730 65
rect 430 15 585 35
rect 655 15 730 35
rect 430 -45 730 15
rect 430 -115 610 -45
rect 630 -115 730 -45
rect 430 -390 730 -115
<< labels >>
rlabel metal1 420 255 420 255 7 VP
port 6 w
rlabel locali 410 -265 410 -265 7 D
port 1 w
rlabel locali 410 -205 410 -205 7 Db
port 2 w
rlabel locali 410 -450 410 -450 7 clk
port 5 w
rlabel metal1 430 -340 430 -340 7 VN
port 7 w
rlabel locali 785 -165 785 -165 3 Q
port 8 e
rlabel locali 785 -265 785 -265 3 Qb
port 9 e
<< end >>
